library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity Aula_12 is
  generic   (
    DATA_WIDTH  : natural :=  32;
    ADDR_WIDTH  : natural :=  32
  );

  port   (
    -- Input ports
    clk     : in  std_logic


  );
end entity;


architecture arch_name of Aula_12 is

	signal flagZero : std_logic;
	signal PC_INC         : std_logic_vector(31 DOWNTO 0);
	signal PC_ROM_INC     : std_logic_vector(31 DOWNTO 0);
	signal PC_ROM         : std_logic_vector(31 DOWNTO 0);
	signal ROM_UC         : std_logic_vector(31 DOWNTO 0);
	signal ULAentradaA_RS : std_logic_vector(31 DOWNTO 0);
	signal ULAentradaB_RT : std_logic_vector(31 DOWNTO 0);
	signal saidaULA       : std_logic_vector(31 DOWNTO 0);
	signal palavraControle_out : std_logic_vector(3 DOWNTO 0);
	
	ALIAS seletor 		           : std_logic_vector(2 DOWNTO 0) IS palavraControle_out(2 DOWNTO 0);
	ALIAS escreveC					  : std_logic IS palavraControle_out(3);
	
	ALIAS entradaA_RS         	  : std_logic_vector (25 DOWNTO 21) IS ROM_UC(25 DOWNTO 21);
	ALIAS entradaB_RT         	  : std_logic_vector (20 DOWNTO 16) IS ROM_UC(20 DOWNTO 16);
	ALIAS entradaC_RD        	  : std_logic_vector (15 DOWNTO 11) IS ROM_UC(15 DOWNTO 11);
	ALIAS opcode            	  : std_logic_vector (31 DOWNTO 26) IS ROM_UC(31 DOWNTO 26);
	ALIAS func            	     : std_logic_vector (5 DOWNTO 0) IS ROM_UC(5 DOWNTO 0);
  
begin

	PC : entity work.registradorGenerico   
						generic map (larguraDados => 32)
						port map (
							DIN => PC_INC, 
							DOUT => PC_ROM_INC, 
							ENABLE => '1', 
							CLK => clk, 
							RST => '0'
						);

	somadorPC : entity work.somaConstante  
						generic map (larguraDados => 32, constante => 4)
						port map( 
							entrada => PC_ROM_INC, 
							saida => PC_INC
						);
							
	ROM_mips: entity work.ROMMIPS
						port map(
							clk => clk,
							Endereco => PC_ROM,
							Dado => ROM_UC
						);
						
	UC: entity work.UnidadeControle
						port map(
							clk => clk,
							opCode => opcode,
							func => func,
							palavraControle => palavraControle_out
						);

	
	bancoRegistrador : entity work.bancoRegistradores   
							 generic map (
								larguraDados => 32, larguraEndBancoRegs => 5 -- 2^5 = 32 posicoes
							)
							 
							 port map ( 
								clk => clk,
								enderecoA => entradaA_RS,
								enderecoB => entradaB_RT,
								enderecoC => entradaC_RD,
								dadoEscritaC => saidaULA,
								escreveC => escreveC,
								saidaA  => ULAentradaA_RS,
								saidaB  => ULAentradaB_RT
								);
	
	
	ULA : entity work.ULA  
							generic map(larguraDados => 32)
							port map (
								entradaA => ULAentradaA_RS, 
								entradaB =>  ULAentradaB_RT,
								saida => saidaULA, 
								seletor => seletor, 
								flagZero => flagZero
								);
							

end architecture;